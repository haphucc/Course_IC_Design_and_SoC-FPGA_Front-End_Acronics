module sqrt_module (
    input wire signed [15:0] delta, // Input delta (16-bit signed)
    output reg [7:0] sqrt_delta      // Square root of delta (8-bit unsigned)
);

    // Lookup table for square roots
    always @(*) begin
        case (delta)
            0: sqrt_delta = 8'd0;
            1: sqrt_delta = 8'd1;
            2, 3: sqrt_delta = 8'd1;
            4: sqrt_delta = 8'd2;
            5, 6, 7, 8: sqrt_delta = 8'd2;
            9: sqrt_delta = 8'd3;
            10, 11, 12, 13, 14, 15: sqrt_delta = 8'd3;
            16: sqrt_delta = 8'd4;
            17, 18, 19, 20, 21, 22, 23, 24: sqrt_delta = 8'd4;
            25: sqrt_delta = 8'd5;
            26, 27, 28, 29, 30, 31, 32, 33, 34, 35: sqrt_delta = 8'd5;
            36: sqrt_delta = 8'd6;
            37, 38, 39, 40, 41, 42, 43, 44, 45, 46, 47, 48: sqrt_delta = 8'd6;
            49: sqrt_delta = 8'd7;
            50, 51, 52, 53, 54, 55, 56, 57, 58, 59, 60, 61, 62, 63, 64: sqrt_delta = 8'd7;
            65, 66, 67, 68, 69, 70, 71, 72, 73, 74, 75, 76, 77, 78, 79, 80: sqrt_delta = 8'd8;
            81: sqrt_delta = 8'd9;
            82, 83, 84, 85, 86, 87, 88, 89, 90, 91, 92, 93, 94, 95, 96, 97, 98, 99, 100: sqrt_delta = 8'd10;
            101, 102, 103, 104, 105, 106, 107, 108, 109, 110, 111, 112, 113, 114, 115, 116, 117, 118, 119, 120, 121: sqrt_delta = 8'd11;
            122, 123, 124, 125, 126, 127, 128, 129, 130, 131, 132, 133, 134, 135, 136, 137, 138, 139, 140, 141, 142, 143, 144: sqrt_delta = 8'd12;
            145, 146, 147, 148, 149, 150, 151, 152, 153, 154, 155, 156, 157, 158, 159, 160, 161, 162, 163, 164, 165, 166, 167, 168, 169: sqrt_delta = 8'd13;
            170, 171, 172, 173, 174, 175, 176, 177, 178, 179, 180, 181, 182, 183, 184, 185, 186, 187, 188, 189, 190, 191, 192, 193, 194, 195, 196: sqrt_delta = 8'd14;
            197, 198, 199, 200, 201, 202, 203, 204, 205, 206, 207, 208, 209, 210, 211, 212, 213, 214, 215, 216, 217, 218, 219, 220, 221, 222, 223, 224, 225: sqrt_delta = 8'd15;
            226, 227, 228, 229, 230, 231, 232, 233, 234, 235, 236, 237, 238, 239, 240, 241, 242, 243, 244, 245, 246, 247, 248, 249, 250, 251, 252, 253, 254, 255, 256: sqrt_delta = 8'd16;
            257, 258, 259, 260, 261, 262, 263, 264, 265, 266, 267, 268, 269, 270, 271, 272, 273, 274, 275, 276, 277, 278, 279, 280, 281, 282, 283, 284, 285, 286, 287, 288, 289: sqrt_delta = 8'd17;
            290, 291, 292, 293, 294, 295, 296, 297, 298, 299, 300, 301, 302, 303, 304, 305, 306, 307, 308, 309, 310, 311, 312, 313, 314, 315, 316, 317, 318, 319, 320, 321, 322, 323, 324: sqrt_delta = 8'd18;
            default: sqrt_delta = 8'd0; // For delta < 0 or > 324
        endcase
    end

endmodule
